-------------------------------------------------------------------------------
--
-- Title       : Fub1
-- Design      : AD7691_VHDL
-- Author      : 
-- Company     : 
--
-------------------------------------------------------------------------------
--
-- File        : C:\My_Designs\MKFP\projekt\AD7691_VHDL\AD7691_VHDL\src\Fub1.vhd
-- Generated   : Thu Jan 26 11:42:49 2017
-- From        : interface description file
-- By          : Itf2Vhdl ver. 1.22
--
-------------------------------------------------------------------------------
--
-- Description : 
--
-------------------------------------------------------------------------------

--{{ Section below this comment is automatically maintained
--   and may be overwritten
--{entity {Fub1} architecture {Fub1}}

library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity Fub1 is
end Fub1;

--}} End of automatically maintained section

architecture Fub1 of Fub1 is
begin

	 -- enter your statements here --

end Fub1;
